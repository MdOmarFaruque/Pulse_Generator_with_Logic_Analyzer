magic
tech sky130A
magscale 1 2
timestamp 1712867557
<< nwell >>
rect 1066 349509 498862 349830
rect 1066 348421 498862 348987
rect 1066 347333 498862 347899
rect 1066 346245 498862 346811
rect 1066 345157 498862 345723
rect 1066 344069 498862 344635
rect 1066 342981 498862 343547
rect 1066 341893 498862 342459
rect 1066 340805 498862 341371
rect 1066 339717 498862 340283
rect 1066 338629 498862 339195
rect 1066 337541 498862 338107
rect 1066 336453 498862 337019
rect 1066 335365 498862 335931
rect 1066 334277 498862 334843
rect 1066 333189 498862 333755
rect 1066 332101 498862 332667
rect 1066 331013 498862 331579
rect 1066 329925 498862 330491
rect 1066 328837 498862 329403
rect 1066 327749 498862 328315
rect 1066 326661 498862 327227
rect 1066 325573 498862 326139
rect 1066 324485 498862 325051
rect 1066 323397 498862 323963
rect 1066 322309 498862 322875
rect 1066 321221 498862 321787
rect 1066 320133 498862 320699
rect 1066 319045 498862 319611
rect 1066 317957 498862 318523
rect 1066 316869 498862 317435
rect 1066 315781 498862 316347
rect 1066 314693 498862 315259
rect 1066 313605 498862 314171
rect 1066 312517 498862 313083
rect 1066 311429 498862 311995
rect 1066 310341 498862 310907
rect 1066 309253 498862 309819
rect 1066 308165 498862 308731
rect 1066 307077 498862 307643
rect 1066 305989 498862 306555
rect 1066 304901 498862 305467
rect 1066 303813 498862 304379
rect 1066 302725 498862 303291
rect 1066 301637 498862 302203
rect 1066 300549 498862 301115
rect 1066 299461 498862 300027
rect 1066 298373 498862 298939
rect 1066 297285 498862 297851
rect 1066 296197 498862 296763
rect 1066 295109 498862 295675
rect 1066 294021 498862 294587
rect 1066 292933 498862 293499
rect 1066 291845 498862 292411
rect 1066 290757 498862 291323
rect 1066 289669 498862 290235
rect 1066 288581 498862 289147
rect 1066 287493 498862 288059
rect 1066 286405 498862 286971
rect 1066 285317 498862 285883
rect 1066 284229 498862 284795
rect 1066 283141 498862 283707
rect 1066 282053 498862 282619
rect 1066 280965 498862 281531
rect 1066 279877 498862 280443
rect 1066 278789 498862 279355
rect 1066 277701 498862 278267
rect 1066 276613 498862 277179
rect 1066 275525 498862 276091
rect 1066 274437 498862 275003
rect 1066 273349 498862 273915
rect 1066 272261 498862 272827
rect 1066 271173 498862 271739
rect 1066 270085 498862 270651
rect 1066 268997 498862 269563
rect 1066 267909 498862 268475
rect 1066 266821 498862 267387
rect 1066 265733 498862 266299
rect 1066 264645 498862 265211
rect 1066 263557 498862 264123
rect 1066 262469 498862 263035
rect 1066 261381 498862 261947
rect 1066 260293 498862 260859
rect 1066 259205 498862 259771
rect 1066 258117 498862 258683
rect 1066 257029 498862 257595
rect 1066 255941 498862 256507
rect 1066 254853 498862 255419
rect 1066 253765 498862 254331
rect 1066 252677 498862 253243
rect 1066 251589 498862 252155
rect 1066 250501 498862 251067
rect 1066 249413 498862 249979
rect 1066 248325 498862 248891
rect 1066 247237 498862 247803
rect 1066 246149 498862 246715
rect 1066 245061 498862 245627
rect 1066 243973 498862 244539
rect 1066 242885 498862 243451
rect 1066 241797 498862 242363
rect 1066 240709 498862 241275
rect 1066 239621 498862 240187
rect 1066 238533 498862 239099
rect 1066 237445 498862 238011
rect 1066 236357 498862 236923
rect 1066 235269 498862 235835
rect 1066 234181 498862 234747
rect 1066 233093 498862 233659
rect 1066 232005 498862 232571
rect 1066 230917 498862 231483
rect 1066 229829 498862 230395
rect 1066 228741 498862 229307
rect 1066 227653 498862 228219
rect 1066 226565 498862 227131
rect 1066 225477 498862 226043
rect 1066 224389 498862 224955
rect 1066 223301 498862 223867
rect 1066 222213 498862 222779
rect 1066 221125 498862 221691
rect 1066 220037 498862 220603
rect 1066 218949 498862 219515
rect 1066 217861 498862 218427
rect 1066 216773 498862 217339
rect 1066 215685 498862 216251
rect 1066 214597 498862 215163
rect 1066 213509 498862 214075
rect 1066 212421 498862 212987
rect 1066 211333 498862 211899
rect 1066 210245 498862 210811
rect 1066 209157 498862 209723
rect 1066 208069 498862 208635
rect 1066 206981 498862 207547
rect 1066 205893 498862 206459
rect 1066 204805 498862 205371
rect 1066 203717 498862 204283
rect 1066 202629 498862 203195
rect 1066 201541 498862 202107
rect 1066 200453 498862 201019
rect 1066 199365 498862 199931
rect 1066 198277 498862 198843
rect 1066 197189 498862 197755
rect 1066 196101 498862 196667
rect 1066 195013 498862 195579
rect 1066 193925 498862 194491
rect 1066 192837 498862 193403
rect 1066 191749 498862 192315
rect 1066 190661 498862 191227
rect 1066 189573 498862 190139
rect 1066 188485 498862 189051
rect 1066 187397 498862 187963
rect 1066 186309 498862 186875
rect 1066 185221 498862 185787
rect 1066 184133 498862 184699
rect 1066 183045 498862 183611
rect 1066 181957 498862 182523
rect 1066 180869 498862 181435
rect 1066 179781 498862 180347
rect 1066 178693 498862 179259
rect 1066 177605 498862 178171
rect 1066 176517 498862 177083
rect 1066 175429 498862 175995
rect 1066 174341 498862 174907
rect 1066 173253 498862 173819
rect 1066 172165 498862 172731
rect 1066 171077 498862 171643
rect 1066 169989 498862 170555
rect 1066 168901 498862 169467
rect 1066 167813 498862 168379
rect 1066 166725 498862 167291
rect 1066 165637 498862 166203
rect 1066 164549 498862 165115
rect 1066 163461 498862 164027
rect 1066 162373 498862 162939
rect 1066 161285 498862 161851
rect 1066 160197 498862 160763
rect 1066 159109 498862 159675
rect 1066 158021 498862 158587
rect 1066 156933 498862 157499
rect 1066 155845 498862 156411
rect 1066 154757 498862 155323
rect 1066 153669 498862 154235
rect 1066 152581 498862 153147
rect 1066 151493 498862 152059
rect 1066 150405 498862 150971
rect 1066 149317 498862 149883
rect 1066 148229 498862 148795
rect 1066 147141 498862 147707
rect 1066 146053 498862 146619
rect 1066 144965 498862 145531
rect 1066 143877 498862 144443
rect 1066 142789 498862 143355
rect 1066 141701 498862 142267
rect 1066 140613 498862 141179
rect 1066 139525 498862 140091
rect 1066 138437 498862 139003
rect 1066 137349 498862 137915
rect 1066 136261 498862 136827
rect 1066 135173 498862 135739
rect 1066 134085 498862 134651
rect 1066 132997 498862 133563
rect 1066 131909 498862 132475
rect 1066 130821 498862 131387
rect 1066 129733 498862 130299
rect 1066 128645 498862 129211
rect 1066 127557 498862 128123
rect 1066 126469 498862 127035
rect 1066 125381 498862 125947
rect 1066 124293 498862 124859
rect 1066 123205 498862 123771
rect 1066 122117 498862 122683
rect 1066 121029 498862 121595
rect 1066 119941 498862 120507
rect 1066 118853 498862 119419
rect 1066 117765 498862 118331
rect 1066 116677 498862 117243
rect 1066 115589 498862 116155
rect 1066 114501 498862 115067
rect 1066 113413 498862 113979
rect 1066 112325 498862 112891
rect 1066 111237 498862 111803
rect 1066 110149 498862 110715
rect 1066 109061 498862 109627
rect 1066 107973 498862 108539
rect 1066 106885 498862 107451
rect 1066 105797 498862 106363
rect 1066 104709 498862 105275
rect 1066 103621 498862 104187
rect 1066 102533 498862 103099
rect 1066 101445 498862 102011
rect 1066 100357 498862 100923
rect 1066 99269 498862 99835
rect 1066 98181 498862 98747
rect 1066 97093 498862 97659
rect 1066 96005 498862 96571
rect 1066 94917 498862 95483
rect 1066 93829 498862 94395
rect 1066 92741 498862 93307
rect 1066 91653 498862 92219
rect 1066 90565 498862 91131
rect 1066 89477 498862 90043
rect 1066 88389 498862 88955
rect 1066 87301 498862 87867
rect 1066 86213 498862 86779
rect 1066 85125 498862 85691
rect 1066 84037 498862 84603
rect 1066 82949 498862 83515
rect 1066 81861 498862 82427
rect 1066 80773 498862 81339
rect 1066 79685 498862 80251
rect 1066 78597 498862 79163
rect 1066 77509 498862 78075
rect 1066 76421 498862 76987
rect 1066 75333 498862 75899
rect 1066 74245 498862 74811
rect 1066 73157 498862 73723
rect 1066 72069 498862 72635
rect 1066 70981 498862 71547
rect 1066 69893 498862 70459
rect 1066 68805 498862 69371
rect 1066 67717 498862 68283
rect 1066 66629 498862 67195
rect 1066 65541 498862 66107
rect 1066 64453 498862 65019
rect 1066 63365 498862 63931
rect 1066 62277 498862 62843
rect 1066 61189 498862 61755
rect 1066 60101 498862 60667
rect 1066 59013 498862 59579
rect 1066 57925 498862 58491
rect 1066 56837 498862 57403
rect 1066 55749 498862 56315
rect 1066 54661 498862 55227
rect 1066 53573 498862 54139
rect 1066 52485 498862 53051
rect 1066 51397 498862 51963
rect 1066 50309 498862 50875
rect 1066 49221 498862 49787
rect 1066 48133 498862 48699
rect 1066 47045 498862 47611
rect 1066 45957 498862 46523
rect 1066 44869 498862 45435
rect 1066 43781 498862 44347
rect 1066 42693 498862 43259
rect 1066 41605 498862 42171
rect 1066 40517 498862 41083
rect 1066 39429 498862 39995
rect 1066 38341 498862 38907
rect 1066 37253 498862 37819
rect 1066 36165 498862 36731
rect 1066 35077 498862 35643
rect 1066 33989 498862 34555
rect 1066 32901 498862 33467
rect 1066 31813 498862 32379
rect 1066 30725 498862 31291
rect 1066 29637 498862 30203
rect 1066 28549 498862 29115
rect 1066 27461 498862 28027
rect 1066 26373 498862 26939
rect 1066 25285 498862 25851
rect 1066 24197 498862 24763
rect 1066 23109 498862 23675
rect 1066 22021 498862 22587
rect 1066 20933 498862 21499
rect 1066 19845 498862 20411
rect 1066 18757 498862 19323
rect 1066 17669 498862 18235
rect 1066 16581 498862 17147
rect 1066 15493 498862 16059
rect 1066 14405 498862 14971
rect 1066 13317 498862 13883
rect 1066 12229 498862 12795
rect 1066 11141 498862 11707
rect 1066 10053 498862 10619
rect 1066 8965 498862 9531
rect 1066 7877 498862 8443
rect 1066 6789 498862 7355
rect 1066 5701 498862 6267
rect 1066 4613 498862 5179
rect 1066 3525 498862 4091
rect 1066 2437 498862 3003
<< obsli1 >>
rect 1104 2159 498824 349809
<< obsm1 >>
rect 1104 1776 498824 349840
<< metal2 >>
rect 17958 0 18014 800
rect 19154 0 19210 800
rect 20350 0 20406 800
rect 21546 0 21602 800
rect 22742 0 22798 800
rect 23938 0 23994 800
rect 25134 0 25190 800
rect 26330 0 26386 800
rect 27526 0 27582 800
rect 28722 0 28778 800
rect 29918 0 29974 800
rect 31114 0 31170 800
rect 32310 0 32366 800
rect 33506 0 33562 800
rect 34702 0 34758 800
rect 35898 0 35954 800
rect 37094 0 37150 800
rect 38290 0 38346 800
rect 39486 0 39542 800
rect 40682 0 40738 800
rect 41878 0 41934 800
rect 43074 0 43130 800
rect 44270 0 44326 800
rect 45466 0 45522 800
rect 46662 0 46718 800
rect 47858 0 47914 800
rect 49054 0 49110 800
rect 50250 0 50306 800
rect 51446 0 51502 800
rect 52642 0 52698 800
rect 53838 0 53894 800
rect 55034 0 55090 800
rect 56230 0 56286 800
rect 57426 0 57482 800
rect 58622 0 58678 800
rect 59818 0 59874 800
rect 61014 0 61070 800
rect 62210 0 62266 800
rect 63406 0 63462 800
rect 64602 0 64658 800
rect 65798 0 65854 800
rect 66994 0 67050 800
rect 68190 0 68246 800
rect 69386 0 69442 800
rect 70582 0 70638 800
rect 71778 0 71834 800
rect 72974 0 73030 800
rect 74170 0 74226 800
rect 75366 0 75422 800
rect 76562 0 76618 800
rect 77758 0 77814 800
rect 78954 0 79010 800
rect 80150 0 80206 800
rect 81346 0 81402 800
rect 82542 0 82598 800
rect 83738 0 83794 800
rect 84934 0 84990 800
rect 86130 0 86186 800
rect 87326 0 87382 800
rect 88522 0 88578 800
rect 89718 0 89774 800
rect 90914 0 90970 800
rect 92110 0 92166 800
rect 93306 0 93362 800
rect 94502 0 94558 800
rect 95698 0 95754 800
rect 96894 0 96950 800
rect 98090 0 98146 800
rect 99286 0 99342 800
rect 100482 0 100538 800
rect 101678 0 101734 800
rect 102874 0 102930 800
rect 104070 0 104126 800
rect 105266 0 105322 800
rect 106462 0 106518 800
rect 107658 0 107714 800
rect 108854 0 108910 800
rect 110050 0 110106 800
rect 111246 0 111302 800
rect 112442 0 112498 800
rect 113638 0 113694 800
rect 114834 0 114890 800
rect 116030 0 116086 800
rect 117226 0 117282 800
rect 118422 0 118478 800
rect 119618 0 119674 800
rect 120814 0 120870 800
rect 122010 0 122066 800
rect 123206 0 123262 800
rect 124402 0 124458 800
rect 125598 0 125654 800
rect 126794 0 126850 800
rect 127990 0 128046 800
rect 129186 0 129242 800
rect 130382 0 130438 800
rect 131578 0 131634 800
rect 132774 0 132830 800
rect 133970 0 134026 800
rect 135166 0 135222 800
rect 136362 0 136418 800
rect 137558 0 137614 800
rect 138754 0 138810 800
rect 139950 0 140006 800
rect 141146 0 141202 800
rect 142342 0 142398 800
rect 143538 0 143594 800
rect 144734 0 144790 800
rect 145930 0 145986 800
rect 147126 0 147182 800
rect 148322 0 148378 800
rect 149518 0 149574 800
rect 150714 0 150770 800
rect 151910 0 151966 800
rect 153106 0 153162 800
rect 154302 0 154358 800
rect 155498 0 155554 800
rect 156694 0 156750 800
rect 157890 0 157946 800
rect 159086 0 159142 800
rect 160282 0 160338 800
rect 161478 0 161534 800
rect 162674 0 162730 800
rect 163870 0 163926 800
rect 165066 0 165122 800
rect 166262 0 166318 800
rect 167458 0 167514 800
rect 168654 0 168710 800
rect 169850 0 169906 800
rect 171046 0 171102 800
rect 172242 0 172298 800
rect 173438 0 173494 800
rect 174634 0 174690 800
rect 175830 0 175886 800
rect 177026 0 177082 800
rect 178222 0 178278 800
rect 179418 0 179474 800
rect 180614 0 180670 800
rect 181810 0 181866 800
rect 183006 0 183062 800
rect 184202 0 184258 800
rect 185398 0 185454 800
rect 186594 0 186650 800
rect 187790 0 187846 800
rect 188986 0 189042 800
rect 190182 0 190238 800
rect 191378 0 191434 800
rect 192574 0 192630 800
rect 193770 0 193826 800
rect 194966 0 195022 800
rect 196162 0 196218 800
rect 197358 0 197414 800
rect 198554 0 198610 800
rect 199750 0 199806 800
rect 200946 0 201002 800
rect 202142 0 202198 800
rect 203338 0 203394 800
rect 204534 0 204590 800
rect 205730 0 205786 800
rect 206926 0 206982 800
rect 208122 0 208178 800
rect 209318 0 209374 800
rect 210514 0 210570 800
rect 211710 0 211766 800
rect 212906 0 212962 800
rect 214102 0 214158 800
rect 215298 0 215354 800
rect 216494 0 216550 800
rect 217690 0 217746 800
rect 218886 0 218942 800
rect 220082 0 220138 800
rect 221278 0 221334 800
rect 222474 0 222530 800
rect 223670 0 223726 800
rect 224866 0 224922 800
rect 226062 0 226118 800
rect 227258 0 227314 800
rect 228454 0 228510 800
rect 229650 0 229706 800
rect 230846 0 230902 800
rect 232042 0 232098 800
rect 233238 0 233294 800
rect 234434 0 234490 800
rect 235630 0 235686 800
rect 236826 0 236882 800
rect 238022 0 238078 800
rect 239218 0 239274 800
rect 240414 0 240470 800
rect 241610 0 241666 800
rect 242806 0 242862 800
rect 244002 0 244058 800
rect 245198 0 245254 800
rect 246394 0 246450 800
rect 247590 0 247646 800
rect 248786 0 248842 800
rect 249982 0 250038 800
rect 251178 0 251234 800
rect 252374 0 252430 800
rect 253570 0 253626 800
rect 254766 0 254822 800
rect 255962 0 256018 800
rect 257158 0 257214 800
rect 258354 0 258410 800
rect 259550 0 259606 800
rect 260746 0 260802 800
rect 261942 0 261998 800
rect 263138 0 263194 800
rect 264334 0 264390 800
rect 265530 0 265586 800
rect 266726 0 266782 800
rect 267922 0 267978 800
rect 269118 0 269174 800
rect 270314 0 270370 800
rect 271510 0 271566 800
rect 272706 0 272762 800
rect 273902 0 273958 800
rect 275098 0 275154 800
rect 276294 0 276350 800
rect 277490 0 277546 800
rect 278686 0 278742 800
rect 279882 0 279938 800
rect 281078 0 281134 800
rect 282274 0 282330 800
rect 283470 0 283526 800
rect 284666 0 284722 800
rect 285862 0 285918 800
rect 287058 0 287114 800
rect 288254 0 288310 800
rect 289450 0 289506 800
rect 290646 0 290702 800
rect 291842 0 291898 800
rect 293038 0 293094 800
rect 294234 0 294290 800
rect 295430 0 295486 800
rect 296626 0 296682 800
rect 297822 0 297878 800
rect 299018 0 299074 800
rect 300214 0 300270 800
rect 301410 0 301466 800
rect 302606 0 302662 800
rect 303802 0 303858 800
rect 304998 0 305054 800
rect 306194 0 306250 800
rect 307390 0 307446 800
rect 308586 0 308642 800
rect 309782 0 309838 800
rect 310978 0 311034 800
rect 312174 0 312230 800
rect 313370 0 313426 800
rect 314566 0 314622 800
rect 315762 0 315818 800
rect 316958 0 317014 800
rect 318154 0 318210 800
rect 319350 0 319406 800
rect 320546 0 320602 800
rect 321742 0 321798 800
rect 322938 0 322994 800
rect 324134 0 324190 800
rect 325330 0 325386 800
rect 326526 0 326582 800
rect 327722 0 327778 800
rect 328918 0 328974 800
rect 330114 0 330170 800
rect 331310 0 331366 800
rect 332506 0 332562 800
rect 333702 0 333758 800
rect 334898 0 334954 800
rect 336094 0 336150 800
rect 337290 0 337346 800
rect 338486 0 338542 800
rect 339682 0 339738 800
rect 340878 0 340934 800
rect 342074 0 342130 800
rect 343270 0 343326 800
rect 344466 0 344522 800
rect 345662 0 345718 800
rect 346858 0 346914 800
rect 348054 0 348110 800
rect 349250 0 349306 800
rect 350446 0 350502 800
rect 351642 0 351698 800
rect 352838 0 352894 800
rect 354034 0 354090 800
rect 355230 0 355286 800
rect 356426 0 356482 800
rect 357622 0 357678 800
rect 358818 0 358874 800
rect 360014 0 360070 800
rect 361210 0 361266 800
rect 362406 0 362462 800
rect 363602 0 363658 800
rect 364798 0 364854 800
rect 365994 0 366050 800
rect 367190 0 367246 800
rect 368386 0 368442 800
rect 369582 0 369638 800
rect 370778 0 370834 800
rect 371974 0 372030 800
rect 373170 0 373226 800
rect 374366 0 374422 800
rect 375562 0 375618 800
rect 376758 0 376814 800
rect 377954 0 378010 800
rect 379150 0 379206 800
rect 380346 0 380402 800
rect 381542 0 381598 800
rect 382738 0 382794 800
rect 383934 0 383990 800
rect 385130 0 385186 800
rect 386326 0 386382 800
rect 387522 0 387578 800
rect 388718 0 388774 800
rect 389914 0 389970 800
rect 391110 0 391166 800
rect 392306 0 392362 800
rect 393502 0 393558 800
rect 394698 0 394754 800
rect 395894 0 395950 800
rect 397090 0 397146 800
rect 398286 0 398342 800
rect 399482 0 399538 800
rect 400678 0 400734 800
rect 401874 0 401930 800
rect 403070 0 403126 800
rect 404266 0 404322 800
rect 405462 0 405518 800
rect 406658 0 406714 800
rect 407854 0 407910 800
rect 409050 0 409106 800
rect 410246 0 410302 800
rect 411442 0 411498 800
rect 412638 0 412694 800
rect 413834 0 413890 800
rect 415030 0 415086 800
rect 416226 0 416282 800
rect 417422 0 417478 800
rect 418618 0 418674 800
rect 419814 0 419870 800
rect 421010 0 421066 800
rect 422206 0 422262 800
rect 423402 0 423458 800
rect 424598 0 424654 800
rect 425794 0 425850 800
rect 426990 0 427046 800
rect 428186 0 428242 800
rect 429382 0 429438 800
rect 430578 0 430634 800
rect 431774 0 431830 800
rect 432970 0 433026 800
rect 434166 0 434222 800
rect 435362 0 435418 800
rect 436558 0 436614 800
rect 437754 0 437810 800
rect 438950 0 439006 800
rect 440146 0 440202 800
rect 441342 0 441398 800
rect 442538 0 442594 800
rect 443734 0 443790 800
rect 444930 0 444986 800
rect 446126 0 446182 800
rect 447322 0 447378 800
rect 448518 0 448574 800
rect 449714 0 449770 800
rect 450910 0 450966 800
rect 452106 0 452162 800
rect 453302 0 453358 800
rect 454498 0 454554 800
rect 455694 0 455750 800
rect 456890 0 456946 800
rect 458086 0 458142 800
rect 459282 0 459338 800
rect 460478 0 460534 800
rect 461674 0 461730 800
rect 462870 0 462926 800
rect 464066 0 464122 800
rect 465262 0 465318 800
rect 466458 0 466514 800
rect 467654 0 467710 800
rect 468850 0 468906 800
rect 470046 0 470102 800
rect 471242 0 471298 800
rect 472438 0 472494 800
rect 473634 0 473690 800
rect 474830 0 474886 800
rect 476026 0 476082 800
rect 477222 0 477278 800
rect 478418 0 478474 800
rect 479614 0 479670 800
rect 480810 0 480866 800
rect 482006 0 482062 800
<< obsm2 >>
rect 4214 856 496042 349829
rect 4214 734 17902 856
rect 18070 734 19098 856
rect 19266 734 20294 856
rect 20462 734 21490 856
rect 21658 734 22686 856
rect 22854 734 23882 856
rect 24050 734 25078 856
rect 25246 734 26274 856
rect 26442 734 27470 856
rect 27638 734 28666 856
rect 28834 734 29862 856
rect 30030 734 31058 856
rect 31226 734 32254 856
rect 32422 734 33450 856
rect 33618 734 34646 856
rect 34814 734 35842 856
rect 36010 734 37038 856
rect 37206 734 38234 856
rect 38402 734 39430 856
rect 39598 734 40626 856
rect 40794 734 41822 856
rect 41990 734 43018 856
rect 43186 734 44214 856
rect 44382 734 45410 856
rect 45578 734 46606 856
rect 46774 734 47802 856
rect 47970 734 48998 856
rect 49166 734 50194 856
rect 50362 734 51390 856
rect 51558 734 52586 856
rect 52754 734 53782 856
rect 53950 734 54978 856
rect 55146 734 56174 856
rect 56342 734 57370 856
rect 57538 734 58566 856
rect 58734 734 59762 856
rect 59930 734 60958 856
rect 61126 734 62154 856
rect 62322 734 63350 856
rect 63518 734 64546 856
rect 64714 734 65742 856
rect 65910 734 66938 856
rect 67106 734 68134 856
rect 68302 734 69330 856
rect 69498 734 70526 856
rect 70694 734 71722 856
rect 71890 734 72918 856
rect 73086 734 74114 856
rect 74282 734 75310 856
rect 75478 734 76506 856
rect 76674 734 77702 856
rect 77870 734 78898 856
rect 79066 734 80094 856
rect 80262 734 81290 856
rect 81458 734 82486 856
rect 82654 734 83682 856
rect 83850 734 84878 856
rect 85046 734 86074 856
rect 86242 734 87270 856
rect 87438 734 88466 856
rect 88634 734 89662 856
rect 89830 734 90858 856
rect 91026 734 92054 856
rect 92222 734 93250 856
rect 93418 734 94446 856
rect 94614 734 95642 856
rect 95810 734 96838 856
rect 97006 734 98034 856
rect 98202 734 99230 856
rect 99398 734 100426 856
rect 100594 734 101622 856
rect 101790 734 102818 856
rect 102986 734 104014 856
rect 104182 734 105210 856
rect 105378 734 106406 856
rect 106574 734 107602 856
rect 107770 734 108798 856
rect 108966 734 109994 856
rect 110162 734 111190 856
rect 111358 734 112386 856
rect 112554 734 113582 856
rect 113750 734 114778 856
rect 114946 734 115974 856
rect 116142 734 117170 856
rect 117338 734 118366 856
rect 118534 734 119562 856
rect 119730 734 120758 856
rect 120926 734 121954 856
rect 122122 734 123150 856
rect 123318 734 124346 856
rect 124514 734 125542 856
rect 125710 734 126738 856
rect 126906 734 127934 856
rect 128102 734 129130 856
rect 129298 734 130326 856
rect 130494 734 131522 856
rect 131690 734 132718 856
rect 132886 734 133914 856
rect 134082 734 135110 856
rect 135278 734 136306 856
rect 136474 734 137502 856
rect 137670 734 138698 856
rect 138866 734 139894 856
rect 140062 734 141090 856
rect 141258 734 142286 856
rect 142454 734 143482 856
rect 143650 734 144678 856
rect 144846 734 145874 856
rect 146042 734 147070 856
rect 147238 734 148266 856
rect 148434 734 149462 856
rect 149630 734 150658 856
rect 150826 734 151854 856
rect 152022 734 153050 856
rect 153218 734 154246 856
rect 154414 734 155442 856
rect 155610 734 156638 856
rect 156806 734 157834 856
rect 158002 734 159030 856
rect 159198 734 160226 856
rect 160394 734 161422 856
rect 161590 734 162618 856
rect 162786 734 163814 856
rect 163982 734 165010 856
rect 165178 734 166206 856
rect 166374 734 167402 856
rect 167570 734 168598 856
rect 168766 734 169794 856
rect 169962 734 170990 856
rect 171158 734 172186 856
rect 172354 734 173382 856
rect 173550 734 174578 856
rect 174746 734 175774 856
rect 175942 734 176970 856
rect 177138 734 178166 856
rect 178334 734 179362 856
rect 179530 734 180558 856
rect 180726 734 181754 856
rect 181922 734 182950 856
rect 183118 734 184146 856
rect 184314 734 185342 856
rect 185510 734 186538 856
rect 186706 734 187734 856
rect 187902 734 188930 856
rect 189098 734 190126 856
rect 190294 734 191322 856
rect 191490 734 192518 856
rect 192686 734 193714 856
rect 193882 734 194910 856
rect 195078 734 196106 856
rect 196274 734 197302 856
rect 197470 734 198498 856
rect 198666 734 199694 856
rect 199862 734 200890 856
rect 201058 734 202086 856
rect 202254 734 203282 856
rect 203450 734 204478 856
rect 204646 734 205674 856
rect 205842 734 206870 856
rect 207038 734 208066 856
rect 208234 734 209262 856
rect 209430 734 210458 856
rect 210626 734 211654 856
rect 211822 734 212850 856
rect 213018 734 214046 856
rect 214214 734 215242 856
rect 215410 734 216438 856
rect 216606 734 217634 856
rect 217802 734 218830 856
rect 218998 734 220026 856
rect 220194 734 221222 856
rect 221390 734 222418 856
rect 222586 734 223614 856
rect 223782 734 224810 856
rect 224978 734 226006 856
rect 226174 734 227202 856
rect 227370 734 228398 856
rect 228566 734 229594 856
rect 229762 734 230790 856
rect 230958 734 231986 856
rect 232154 734 233182 856
rect 233350 734 234378 856
rect 234546 734 235574 856
rect 235742 734 236770 856
rect 236938 734 237966 856
rect 238134 734 239162 856
rect 239330 734 240358 856
rect 240526 734 241554 856
rect 241722 734 242750 856
rect 242918 734 243946 856
rect 244114 734 245142 856
rect 245310 734 246338 856
rect 246506 734 247534 856
rect 247702 734 248730 856
rect 248898 734 249926 856
rect 250094 734 251122 856
rect 251290 734 252318 856
rect 252486 734 253514 856
rect 253682 734 254710 856
rect 254878 734 255906 856
rect 256074 734 257102 856
rect 257270 734 258298 856
rect 258466 734 259494 856
rect 259662 734 260690 856
rect 260858 734 261886 856
rect 262054 734 263082 856
rect 263250 734 264278 856
rect 264446 734 265474 856
rect 265642 734 266670 856
rect 266838 734 267866 856
rect 268034 734 269062 856
rect 269230 734 270258 856
rect 270426 734 271454 856
rect 271622 734 272650 856
rect 272818 734 273846 856
rect 274014 734 275042 856
rect 275210 734 276238 856
rect 276406 734 277434 856
rect 277602 734 278630 856
rect 278798 734 279826 856
rect 279994 734 281022 856
rect 281190 734 282218 856
rect 282386 734 283414 856
rect 283582 734 284610 856
rect 284778 734 285806 856
rect 285974 734 287002 856
rect 287170 734 288198 856
rect 288366 734 289394 856
rect 289562 734 290590 856
rect 290758 734 291786 856
rect 291954 734 292982 856
rect 293150 734 294178 856
rect 294346 734 295374 856
rect 295542 734 296570 856
rect 296738 734 297766 856
rect 297934 734 298962 856
rect 299130 734 300158 856
rect 300326 734 301354 856
rect 301522 734 302550 856
rect 302718 734 303746 856
rect 303914 734 304942 856
rect 305110 734 306138 856
rect 306306 734 307334 856
rect 307502 734 308530 856
rect 308698 734 309726 856
rect 309894 734 310922 856
rect 311090 734 312118 856
rect 312286 734 313314 856
rect 313482 734 314510 856
rect 314678 734 315706 856
rect 315874 734 316902 856
rect 317070 734 318098 856
rect 318266 734 319294 856
rect 319462 734 320490 856
rect 320658 734 321686 856
rect 321854 734 322882 856
rect 323050 734 324078 856
rect 324246 734 325274 856
rect 325442 734 326470 856
rect 326638 734 327666 856
rect 327834 734 328862 856
rect 329030 734 330058 856
rect 330226 734 331254 856
rect 331422 734 332450 856
rect 332618 734 333646 856
rect 333814 734 334842 856
rect 335010 734 336038 856
rect 336206 734 337234 856
rect 337402 734 338430 856
rect 338598 734 339626 856
rect 339794 734 340822 856
rect 340990 734 342018 856
rect 342186 734 343214 856
rect 343382 734 344410 856
rect 344578 734 345606 856
rect 345774 734 346802 856
rect 346970 734 347998 856
rect 348166 734 349194 856
rect 349362 734 350390 856
rect 350558 734 351586 856
rect 351754 734 352782 856
rect 352950 734 353978 856
rect 354146 734 355174 856
rect 355342 734 356370 856
rect 356538 734 357566 856
rect 357734 734 358762 856
rect 358930 734 359958 856
rect 360126 734 361154 856
rect 361322 734 362350 856
rect 362518 734 363546 856
rect 363714 734 364742 856
rect 364910 734 365938 856
rect 366106 734 367134 856
rect 367302 734 368330 856
rect 368498 734 369526 856
rect 369694 734 370722 856
rect 370890 734 371918 856
rect 372086 734 373114 856
rect 373282 734 374310 856
rect 374478 734 375506 856
rect 375674 734 376702 856
rect 376870 734 377898 856
rect 378066 734 379094 856
rect 379262 734 380290 856
rect 380458 734 381486 856
rect 381654 734 382682 856
rect 382850 734 383878 856
rect 384046 734 385074 856
rect 385242 734 386270 856
rect 386438 734 387466 856
rect 387634 734 388662 856
rect 388830 734 389858 856
rect 390026 734 391054 856
rect 391222 734 392250 856
rect 392418 734 393446 856
rect 393614 734 394642 856
rect 394810 734 395838 856
rect 396006 734 397034 856
rect 397202 734 398230 856
rect 398398 734 399426 856
rect 399594 734 400622 856
rect 400790 734 401818 856
rect 401986 734 403014 856
rect 403182 734 404210 856
rect 404378 734 405406 856
rect 405574 734 406602 856
rect 406770 734 407798 856
rect 407966 734 408994 856
rect 409162 734 410190 856
rect 410358 734 411386 856
rect 411554 734 412582 856
rect 412750 734 413778 856
rect 413946 734 414974 856
rect 415142 734 416170 856
rect 416338 734 417366 856
rect 417534 734 418562 856
rect 418730 734 419758 856
rect 419926 734 420954 856
rect 421122 734 422150 856
rect 422318 734 423346 856
rect 423514 734 424542 856
rect 424710 734 425738 856
rect 425906 734 426934 856
rect 427102 734 428130 856
rect 428298 734 429326 856
rect 429494 734 430522 856
rect 430690 734 431718 856
rect 431886 734 432914 856
rect 433082 734 434110 856
rect 434278 734 435306 856
rect 435474 734 436502 856
rect 436670 734 437698 856
rect 437866 734 438894 856
rect 439062 734 440090 856
rect 440258 734 441286 856
rect 441454 734 442482 856
rect 442650 734 443678 856
rect 443846 734 444874 856
rect 445042 734 446070 856
rect 446238 734 447266 856
rect 447434 734 448462 856
rect 448630 734 449658 856
rect 449826 734 450854 856
rect 451022 734 452050 856
rect 452218 734 453246 856
rect 453414 734 454442 856
rect 454610 734 455638 856
rect 455806 734 456834 856
rect 457002 734 458030 856
rect 458198 734 459226 856
rect 459394 734 460422 856
rect 460590 734 461618 856
rect 461786 734 462814 856
rect 462982 734 464010 856
rect 464178 734 465206 856
rect 465374 734 466402 856
rect 466570 734 467598 856
rect 467766 734 468794 856
rect 468962 734 469990 856
rect 470158 734 471186 856
rect 471354 734 472382 856
rect 472550 734 473578 856
rect 473746 734 474774 856
rect 474942 734 475970 856
rect 476138 734 477166 856
rect 477334 734 478362 856
rect 478530 734 479558 856
rect 479726 734 480754 856
rect 480922 734 481950 856
rect 482118 734 496042 856
<< obsm3 >>
rect 4210 2143 496046 349825
<< metal4 >>
rect 4208 2128 4528 349840
rect 11888 2128 12208 349840
rect 19568 2128 19888 349840
rect 27248 2128 27568 349840
rect 34928 2128 35248 349840
rect 42608 2128 42928 349840
rect 50288 2128 50608 349840
rect 57968 2128 58288 349840
rect 65648 2128 65968 349840
rect 73328 2128 73648 349840
rect 81008 2128 81328 349840
rect 88688 2128 89008 349840
rect 96368 2128 96688 349840
rect 104048 2128 104368 349840
rect 111728 2128 112048 349840
rect 119408 2128 119728 349840
rect 127088 2128 127408 349840
rect 134768 2128 135088 349840
rect 142448 2128 142768 349840
rect 150128 2128 150448 349840
rect 157808 2128 158128 349840
rect 165488 2128 165808 349840
rect 173168 2128 173488 349840
rect 180848 2128 181168 349840
rect 188528 2128 188848 349840
rect 196208 2128 196528 349840
rect 203888 2128 204208 349840
rect 211568 2128 211888 349840
rect 219248 2128 219568 349840
rect 226928 2128 227248 349840
rect 234608 2128 234928 349840
rect 242288 2128 242608 349840
rect 249968 2128 250288 349840
rect 257648 2128 257968 349840
rect 265328 2128 265648 349840
rect 273008 2128 273328 349840
rect 280688 2128 281008 349840
rect 288368 2128 288688 349840
rect 296048 2128 296368 349840
rect 303728 2128 304048 349840
rect 311408 2128 311728 349840
rect 319088 2128 319408 349840
rect 326768 2128 327088 349840
rect 334448 2128 334768 349840
rect 342128 2128 342448 349840
rect 349808 2128 350128 349840
rect 357488 2128 357808 349840
rect 365168 2128 365488 349840
rect 372848 2128 373168 349840
rect 380528 2128 380848 349840
rect 388208 2128 388528 349840
rect 395888 2128 396208 349840
rect 403568 2128 403888 349840
rect 411248 2128 411568 349840
rect 418928 2128 419248 349840
rect 426608 2128 426928 349840
rect 434288 2128 434608 349840
rect 441968 2128 442288 349840
rect 449648 2128 449968 349840
rect 457328 2128 457648 349840
rect 465008 2128 465328 349840
rect 472688 2128 473008 349840
rect 480368 2128 480688 349840
rect 488048 2128 488368 349840
rect 495728 2128 496048 349840
<< labels >>
rlabel metal2 s 482006 0 482062 800 6 analog_io2
port 1 nsew signal output
rlabel metal2 s 22742 0 22798 800 6 la_data_in[0]
port 2 nsew signal input
rlabel metal2 s 381542 0 381598 800 6 la_data_in[100]
port 3 nsew signal input
rlabel metal2 s 385130 0 385186 800 6 la_data_in[101]
port 4 nsew signal input
rlabel metal2 s 388718 0 388774 800 6 la_data_in[102]
port 5 nsew signal input
rlabel metal2 s 392306 0 392362 800 6 la_data_in[103]
port 6 nsew signal input
rlabel metal2 s 395894 0 395950 800 6 la_data_in[104]
port 7 nsew signal input
rlabel metal2 s 399482 0 399538 800 6 la_data_in[105]
port 8 nsew signal input
rlabel metal2 s 403070 0 403126 800 6 la_data_in[106]
port 9 nsew signal input
rlabel metal2 s 406658 0 406714 800 6 la_data_in[107]
port 10 nsew signal input
rlabel metal2 s 410246 0 410302 800 6 la_data_in[108]
port 11 nsew signal input
rlabel metal2 s 413834 0 413890 800 6 la_data_in[109]
port 12 nsew signal input
rlabel metal2 s 58622 0 58678 800 6 la_data_in[10]
port 13 nsew signal input
rlabel metal2 s 417422 0 417478 800 6 la_data_in[110]
port 14 nsew signal input
rlabel metal2 s 421010 0 421066 800 6 la_data_in[111]
port 15 nsew signal input
rlabel metal2 s 424598 0 424654 800 6 la_data_in[112]
port 16 nsew signal input
rlabel metal2 s 428186 0 428242 800 6 la_data_in[113]
port 17 nsew signal input
rlabel metal2 s 431774 0 431830 800 6 la_data_in[114]
port 18 nsew signal input
rlabel metal2 s 435362 0 435418 800 6 la_data_in[115]
port 19 nsew signal input
rlabel metal2 s 438950 0 439006 800 6 la_data_in[116]
port 20 nsew signal input
rlabel metal2 s 442538 0 442594 800 6 la_data_in[117]
port 21 nsew signal input
rlabel metal2 s 446126 0 446182 800 6 la_data_in[118]
port 22 nsew signal input
rlabel metal2 s 449714 0 449770 800 6 la_data_in[119]
port 23 nsew signal input
rlabel metal2 s 62210 0 62266 800 6 la_data_in[11]
port 24 nsew signal input
rlabel metal2 s 453302 0 453358 800 6 la_data_in[120]
port 25 nsew signal input
rlabel metal2 s 456890 0 456946 800 6 la_data_in[121]
port 26 nsew signal input
rlabel metal2 s 460478 0 460534 800 6 la_data_in[122]
port 27 nsew signal input
rlabel metal2 s 464066 0 464122 800 6 la_data_in[123]
port 28 nsew signal input
rlabel metal2 s 467654 0 467710 800 6 la_data_in[124]
port 29 nsew signal input
rlabel metal2 s 471242 0 471298 800 6 la_data_in[125]
port 30 nsew signal input
rlabel metal2 s 474830 0 474886 800 6 la_data_in[126]
port 31 nsew signal input
rlabel metal2 s 478418 0 478474 800 6 la_data_in[127]
port 32 nsew signal input
rlabel metal2 s 65798 0 65854 800 6 la_data_in[12]
port 33 nsew signal input
rlabel metal2 s 69386 0 69442 800 6 la_data_in[13]
port 34 nsew signal input
rlabel metal2 s 72974 0 73030 800 6 la_data_in[14]
port 35 nsew signal input
rlabel metal2 s 76562 0 76618 800 6 la_data_in[15]
port 36 nsew signal input
rlabel metal2 s 80150 0 80206 800 6 la_data_in[16]
port 37 nsew signal input
rlabel metal2 s 83738 0 83794 800 6 la_data_in[17]
port 38 nsew signal input
rlabel metal2 s 87326 0 87382 800 6 la_data_in[18]
port 39 nsew signal input
rlabel metal2 s 90914 0 90970 800 6 la_data_in[19]
port 40 nsew signal input
rlabel metal2 s 26330 0 26386 800 6 la_data_in[1]
port 41 nsew signal input
rlabel metal2 s 94502 0 94558 800 6 la_data_in[20]
port 42 nsew signal input
rlabel metal2 s 98090 0 98146 800 6 la_data_in[21]
port 43 nsew signal input
rlabel metal2 s 101678 0 101734 800 6 la_data_in[22]
port 44 nsew signal input
rlabel metal2 s 105266 0 105322 800 6 la_data_in[23]
port 45 nsew signal input
rlabel metal2 s 108854 0 108910 800 6 la_data_in[24]
port 46 nsew signal input
rlabel metal2 s 112442 0 112498 800 6 la_data_in[25]
port 47 nsew signal input
rlabel metal2 s 116030 0 116086 800 6 la_data_in[26]
port 48 nsew signal input
rlabel metal2 s 119618 0 119674 800 6 la_data_in[27]
port 49 nsew signal input
rlabel metal2 s 123206 0 123262 800 6 la_data_in[28]
port 50 nsew signal input
rlabel metal2 s 126794 0 126850 800 6 la_data_in[29]
port 51 nsew signal input
rlabel metal2 s 29918 0 29974 800 6 la_data_in[2]
port 52 nsew signal input
rlabel metal2 s 130382 0 130438 800 6 la_data_in[30]
port 53 nsew signal input
rlabel metal2 s 133970 0 134026 800 6 la_data_in[31]
port 54 nsew signal input
rlabel metal2 s 137558 0 137614 800 6 la_data_in[32]
port 55 nsew signal input
rlabel metal2 s 141146 0 141202 800 6 la_data_in[33]
port 56 nsew signal input
rlabel metal2 s 144734 0 144790 800 6 la_data_in[34]
port 57 nsew signal input
rlabel metal2 s 148322 0 148378 800 6 la_data_in[35]
port 58 nsew signal input
rlabel metal2 s 151910 0 151966 800 6 la_data_in[36]
port 59 nsew signal input
rlabel metal2 s 155498 0 155554 800 6 la_data_in[37]
port 60 nsew signal input
rlabel metal2 s 159086 0 159142 800 6 la_data_in[38]
port 61 nsew signal input
rlabel metal2 s 162674 0 162730 800 6 la_data_in[39]
port 62 nsew signal input
rlabel metal2 s 33506 0 33562 800 6 la_data_in[3]
port 63 nsew signal input
rlabel metal2 s 166262 0 166318 800 6 la_data_in[40]
port 64 nsew signal input
rlabel metal2 s 169850 0 169906 800 6 la_data_in[41]
port 65 nsew signal input
rlabel metal2 s 173438 0 173494 800 6 la_data_in[42]
port 66 nsew signal input
rlabel metal2 s 177026 0 177082 800 6 la_data_in[43]
port 67 nsew signal input
rlabel metal2 s 180614 0 180670 800 6 la_data_in[44]
port 68 nsew signal input
rlabel metal2 s 184202 0 184258 800 6 la_data_in[45]
port 69 nsew signal input
rlabel metal2 s 187790 0 187846 800 6 la_data_in[46]
port 70 nsew signal input
rlabel metal2 s 191378 0 191434 800 6 la_data_in[47]
port 71 nsew signal input
rlabel metal2 s 194966 0 195022 800 6 la_data_in[48]
port 72 nsew signal input
rlabel metal2 s 198554 0 198610 800 6 la_data_in[49]
port 73 nsew signal input
rlabel metal2 s 37094 0 37150 800 6 la_data_in[4]
port 74 nsew signal input
rlabel metal2 s 202142 0 202198 800 6 la_data_in[50]
port 75 nsew signal input
rlabel metal2 s 205730 0 205786 800 6 la_data_in[51]
port 76 nsew signal input
rlabel metal2 s 209318 0 209374 800 6 la_data_in[52]
port 77 nsew signal input
rlabel metal2 s 212906 0 212962 800 6 la_data_in[53]
port 78 nsew signal input
rlabel metal2 s 216494 0 216550 800 6 la_data_in[54]
port 79 nsew signal input
rlabel metal2 s 220082 0 220138 800 6 la_data_in[55]
port 80 nsew signal input
rlabel metal2 s 223670 0 223726 800 6 la_data_in[56]
port 81 nsew signal input
rlabel metal2 s 227258 0 227314 800 6 la_data_in[57]
port 82 nsew signal input
rlabel metal2 s 230846 0 230902 800 6 la_data_in[58]
port 83 nsew signal input
rlabel metal2 s 234434 0 234490 800 6 la_data_in[59]
port 84 nsew signal input
rlabel metal2 s 40682 0 40738 800 6 la_data_in[5]
port 85 nsew signal input
rlabel metal2 s 238022 0 238078 800 6 la_data_in[60]
port 86 nsew signal input
rlabel metal2 s 241610 0 241666 800 6 la_data_in[61]
port 87 nsew signal input
rlabel metal2 s 245198 0 245254 800 6 la_data_in[62]
port 88 nsew signal input
rlabel metal2 s 248786 0 248842 800 6 la_data_in[63]
port 89 nsew signal input
rlabel metal2 s 252374 0 252430 800 6 la_data_in[64]
port 90 nsew signal input
rlabel metal2 s 255962 0 256018 800 6 la_data_in[65]
port 91 nsew signal input
rlabel metal2 s 259550 0 259606 800 6 la_data_in[66]
port 92 nsew signal input
rlabel metal2 s 263138 0 263194 800 6 la_data_in[67]
port 93 nsew signal input
rlabel metal2 s 266726 0 266782 800 6 la_data_in[68]
port 94 nsew signal input
rlabel metal2 s 270314 0 270370 800 6 la_data_in[69]
port 95 nsew signal input
rlabel metal2 s 44270 0 44326 800 6 la_data_in[6]
port 96 nsew signal input
rlabel metal2 s 273902 0 273958 800 6 la_data_in[70]
port 97 nsew signal input
rlabel metal2 s 277490 0 277546 800 6 la_data_in[71]
port 98 nsew signal input
rlabel metal2 s 281078 0 281134 800 6 la_data_in[72]
port 99 nsew signal input
rlabel metal2 s 284666 0 284722 800 6 la_data_in[73]
port 100 nsew signal input
rlabel metal2 s 288254 0 288310 800 6 la_data_in[74]
port 101 nsew signal input
rlabel metal2 s 291842 0 291898 800 6 la_data_in[75]
port 102 nsew signal input
rlabel metal2 s 295430 0 295486 800 6 la_data_in[76]
port 103 nsew signal input
rlabel metal2 s 299018 0 299074 800 6 la_data_in[77]
port 104 nsew signal input
rlabel metal2 s 302606 0 302662 800 6 la_data_in[78]
port 105 nsew signal input
rlabel metal2 s 306194 0 306250 800 6 la_data_in[79]
port 106 nsew signal input
rlabel metal2 s 47858 0 47914 800 6 la_data_in[7]
port 107 nsew signal input
rlabel metal2 s 309782 0 309838 800 6 la_data_in[80]
port 108 nsew signal input
rlabel metal2 s 313370 0 313426 800 6 la_data_in[81]
port 109 nsew signal input
rlabel metal2 s 316958 0 317014 800 6 la_data_in[82]
port 110 nsew signal input
rlabel metal2 s 320546 0 320602 800 6 la_data_in[83]
port 111 nsew signal input
rlabel metal2 s 324134 0 324190 800 6 la_data_in[84]
port 112 nsew signal input
rlabel metal2 s 327722 0 327778 800 6 la_data_in[85]
port 113 nsew signal input
rlabel metal2 s 331310 0 331366 800 6 la_data_in[86]
port 114 nsew signal input
rlabel metal2 s 334898 0 334954 800 6 la_data_in[87]
port 115 nsew signal input
rlabel metal2 s 338486 0 338542 800 6 la_data_in[88]
port 116 nsew signal input
rlabel metal2 s 342074 0 342130 800 6 la_data_in[89]
port 117 nsew signal input
rlabel metal2 s 51446 0 51502 800 6 la_data_in[8]
port 118 nsew signal input
rlabel metal2 s 345662 0 345718 800 6 la_data_in[90]
port 119 nsew signal input
rlabel metal2 s 349250 0 349306 800 6 la_data_in[91]
port 120 nsew signal input
rlabel metal2 s 352838 0 352894 800 6 la_data_in[92]
port 121 nsew signal input
rlabel metal2 s 356426 0 356482 800 6 la_data_in[93]
port 122 nsew signal input
rlabel metal2 s 360014 0 360070 800 6 la_data_in[94]
port 123 nsew signal input
rlabel metal2 s 363602 0 363658 800 6 la_data_in[95]
port 124 nsew signal input
rlabel metal2 s 367190 0 367246 800 6 la_data_in[96]
port 125 nsew signal input
rlabel metal2 s 370778 0 370834 800 6 la_data_in[97]
port 126 nsew signal input
rlabel metal2 s 374366 0 374422 800 6 la_data_in[98]
port 127 nsew signal input
rlabel metal2 s 377954 0 378010 800 6 la_data_in[99]
port 128 nsew signal input
rlabel metal2 s 55034 0 55090 800 6 la_data_in[9]
port 129 nsew signal input
rlabel metal2 s 23938 0 23994 800 6 la_data_out[0]
port 130 nsew signal output
rlabel metal2 s 382738 0 382794 800 6 la_data_out[100]
port 131 nsew signal output
rlabel metal2 s 386326 0 386382 800 6 la_data_out[101]
port 132 nsew signal output
rlabel metal2 s 389914 0 389970 800 6 la_data_out[102]
port 133 nsew signal output
rlabel metal2 s 393502 0 393558 800 6 la_data_out[103]
port 134 nsew signal output
rlabel metal2 s 397090 0 397146 800 6 la_data_out[104]
port 135 nsew signal output
rlabel metal2 s 400678 0 400734 800 6 la_data_out[105]
port 136 nsew signal output
rlabel metal2 s 404266 0 404322 800 6 la_data_out[106]
port 137 nsew signal output
rlabel metal2 s 407854 0 407910 800 6 la_data_out[107]
port 138 nsew signal output
rlabel metal2 s 411442 0 411498 800 6 la_data_out[108]
port 139 nsew signal output
rlabel metal2 s 415030 0 415086 800 6 la_data_out[109]
port 140 nsew signal output
rlabel metal2 s 59818 0 59874 800 6 la_data_out[10]
port 141 nsew signal output
rlabel metal2 s 418618 0 418674 800 6 la_data_out[110]
port 142 nsew signal output
rlabel metal2 s 422206 0 422262 800 6 la_data_out[111]
port 143 nsew signal output
rlabel metal2 s 425794 0 425850 800 6 la_data_out[112]
port 144 nsew signal output
rlabel metal2 s 429382 0 429438 800 6 la_data_out[113]
port 145 nsew signal output
rlabel metal2 s 432970 0 433026 800 6 la_data_out[114]
port 146 nsew signal output
rlabel metal2 s 436558 0 436614 800 6 la_data_out[115]
port 147 nsew signal output
rlabel metal2 s 440146 0 440202 800 6 la_data_out[116]
port 148 nsew signal output
rlabel metal2 s 443734 0 443790 800 6 la_data_out[117]
port 149 nsew signal output
rlabel metal2 s 447322 0 447378 800 6 la_data_out[118]
port 150 nsew signal output
rlabel metal2 s 450910 0 450966 800 6 la_data_out[119]
port 151 nsew signal output
rlabel metal2 s 63406 0 63462 800 6 la_data_out[11]
port 152 nsew signal output
rlabel metal2 s 454498 0 454554 800 6 la_data_out[120]
port 153 nsew signal output
rlabel metal2 s 458086 0 458142 800 6 la_data_out[121]
port 154 nsew signal output
rlabel metal2 s 461674 0 461730 800 6 la_data_out[122]
port 155 nsew signal output
rlabel metal2 s 465262 0 465318 800 6 la_data_out[123]
port 156 nsew signal output
rlabel metal2 s 468850 0 468906 800 6 la_data_out[124]
port 157 nsew signal output
rlabel metal2 s 472438 0 472494 800 6 la_data_out[125]
port 158 nsew signal output
rlabel metal2 s 476026 0 476082 800 6 la_data_out[126]
port 159 nsew signal output
rlabel metal2 s 479614 0 479670 800 6 la_data_out[127]
port 160 nsew signal output
rlabel metal2 s 66994 0 67050 800 6 la_data_out[12]
port 161 nsew signal output
rlabel metal2 s 70582 0 70638 800 6 la_data_out[13]
port 162 nsew signal output
rlabel metal2 s 74170 0 74226 800 6 la_data_out[14]
port 163 nsew signal output
rlabel metal2 s 77758 0 77814 800 6 la_data_out[15]
port 164 nsew signal output
rlabel metal2 s 81346 0 81402 800 6 la_data_out[16]
port 165 nsew signal output
rlabel metal2 s 84934 0 84990 800 6 la_data_out[17]
port 166 nsew signal output
rlabel metal2 s 88522 0 88578 800 6 la_data_out[18]
port 167 nsew signal output
rlabel metal2 s 92110 0 92166 800 6 la_data_out[19]
port 168 nsew signal output
rlabel metal2 s 27526 0 27582 800 6 la_data_out[1]
port 169 nsew signal output
rlabel metal2 s 95698 0 95754 800 6 la_data_out[20]
port 170 nsew signal output
rlabel metal2 s 99286 0 99342 800 6 la_data_out[21]
port 171 nsew signal output
rlabel metal2 s 102874 0 102930 800 6 la_data_out[22]
port 172 nsew signal output
rlabel metal2 s 106462 0 106518 800 6 la_data_out[23]
port 173 nsew signal output
rlabel metal2 s 110050 0 110106 800 6 la_data_out[24]
port 174 nsew signal output
rlabel metal2 s 113638 0 113694 800 6 la_data_out[25]
port 175 nsew signal output
rlabel metal2 s 117226 0 117282 800 6 la_data_out[26]
port 176 nsew signal output
rlabel metal2 s 120814 0 120870 800 6 la_data_out[27]
port 177 nsew signal output
rlabel metal2 s 124402 0 124458 800 6 la_data_out[28]
port 178 nsew signal output
rlabel metal2 s 127990 0 128046 800 6 la_data_out[29]
port 179 nsew signal output
rlabel metal2 s 31114 0 31170 800 6 la_data_out[2]
port 180 nsew signal output
rlabel metal2 s 131578 0 131634 800 6 la_data_out[30]
port 181 nsew signal output
rlabel metal2 s 135166 0 135222 800 6 la_data_out[31]
port 182 nsew signal output
rlabel metal2 s 138754 0 138810 800 6 la_data_out[32]
port 183 nsew signal output
rlabel metal2 s 142342 0 142398 800 6 la_data_out[33]
port 184 nsew signal output
rlabel metal2 s 145930 0 145986 800 6 la_data_out[34]
port 185 nsew signal output
rlabel metal2 s 149518 0 149574 800 6 la_data_out[35]
port 186 nsew signal output
rlabel metal2 s 153106 0 153162 800 6 la_data_out[36]
port 187 nsew signal output
rlabel metal2 s 156694 0 156750 800 6 la_data_out[37]
port 188 nsew signal output
rlabel metal2 s 160282 0 160338 800 6 la_data_out[38]
port 189 nsew signal output
rlabel metal2 s 163870 0 163926 800 6 la_data_out[39]
port 190 nsew signal output
rlabel metal2 s 34702 0 34758 800 6 la_data_out[3]
port 191 nsew signal output
rlabel metal2 s 167458 0 167514 800 6 la_data_out[40]
port 192 nsew signal output
rlabel metal2 s 171046 0 171102 800 6 la_data_out[41]
port 193 nsew signal output
rlabel metal2 s 174634 0 174690 800 6 la_data_out[42]
port 194 nsew signal output
rlabel metal2 s 178222 0 178278 800 6 la_data_out[43]
port 195 nsew signal output
rlabel metal2 s 181810 0 181866 800 6 la_data_out[44]
port 196 nsew signal output
rlabel metal2 s 185398 0 185454 800 6 la_data_out[45]
port 197 nsew signal output
rlabel metal2 s 188986 0 189042 800 6 la_data_out[46]
port 198 nsew signal output
rlabel metal2 s 192574 0 192630 800 6 la_data_out[47]
port 199 nsew signal output
rlabel metal2 s 196162 0 196218 800 6 la_data_out[48]
port 200 nsew signal output
rlabel metal2 s 199750 0 199806 800 6 la_data_out[49]
port 201 nsew signal output
rlabel metal2 s 38290 0 38346 800 6 la_data_out[4]
port 202 nsew signal output
rlabel metal2 s 203338 0 203394 800 6 la_data_out[50]
port 203 nsew signal output
rlabel metal2 s 206926 0 206982 800 6 la_data_out[51]
port 204 nsew signal output
rlabel metal2 s 210514 0 210570 800 6 la_data_out[52]
port 205 nsew signal output
rlabel metal2 s 214102 0 214158 800 6 la_data_out[53]
port 206 nsew signal output
rlabel metal2 s 217690 0 217746 800 6 la_data_out[54]
port 207 nsew signal output
rlabel metal2 s 221278 0 221334 800 6 la_data_out[55]
port 208 nsew signal output
rlabel metal2 s 224866 0 224922 800 6 la_data_out[56]
port 209 nsew signal output
rlabel metal2 s 228454 0 228510 800 6 la_data_out[57]
port 210 nsew signal output
rlabel metal2 s 232042 0 232098 800 6 la_data_out[58]
port 211 nsew signal output
rlabel metal2 s 235630 0 235686 800 6 la_data_out[59]
port 212 nsew signal output
rlabel metal2 s 41878 0 41934 800 6 la_data_out[5]
port 213 nsew signal output
rlabel metal2 s 239218 0 239274 800 6 la_data_out[60]
port 214 nsew signal output
rlabel metal2 s 242806 0 242862 800 6 la_data_out[61]
port 215 nsew signal output
rlabel metal2 s 246394 0 246450 800 6 la_data_out[62]
port 216 nsew signal output
rlabel metal2 s 249982 0 250038 800 6 la_data_out[63]
port 217 nsew signal output
rlabel metal2 s 253570 0 253626 800 6 la_data_out[64]
port 218 nsew signal output
rlabel metal2 s 257158 0 257214 800 6 la_data_out[65]
port 219 nsew signal output
rlabel metal2 s 260746 0 260802 800 6 la_data_out[66]
port 220 nsew signal output
rlabel metal2 s 264334 0 264390 800 6 la_data_out[67]
port 221 nsew signal output
rlabel metal2 s 267922 0 267978 800 6 la_data_out[68]
port 222 nsew signal output
rlabel metal2 s 271510 0 271566 800 6 la_data_out[69]
port 223 nsew signal output
rlabel metal2 s 45466 0 45522 800 6 la_data_out[6]
port 224 nsew signal output
rlabel metal2 s 275098 0 275154 800 6 la_data_out[70]
port 225 nsew signal output
rlabel metal2 s 278686 0 278742 800 6 la_data_out[71]
port 226 nsew signal output
rlabel metal2 s 282274 0 282330 800 6 la_data_out[72]
port 227 nsew signal output
rlabel metal2 s 285862 0 285918 800 6 la_data_out[73]
port 228 nsew signal output
rlabel metal2 s 289450 0 289506 800 6 la_data_out[74]
port 229 nsew signal output
rlabel metal2 s 293038 0 293094 800 6 la_data_out[75]
port 230 nsew signal output
rlabel metal2 s 296626 0 296682 800 6 la_data_out[76]
port 231 nsew signal output
rlabel metal2 s 300214 0 300270 800 6 la_data_out[77]
port 232 nsew signal output
rlabel metal2 s 303802 0 303858 800 6 la_data_out[78]
port 233 nsew signal output
rlabel metal2 s 307390 0 307446 800 6 la_data_out[79]
port 234 nsew signal output
rlabel metal2 s 49054 0 49110 800 6 la_data_out[7]
port 235 nsew signal output
rlabel metal2 s 310978 0 311034 800 6 la_data_out[80]
port 236 nsew signal output
rlabel metal2 s 314566 0 314622 800 6 la_data_out[81]
port 237 nsew signal output
rlabel metal2 s 318154 0 318210 800 6 la_data_out[82]
port 238 nsew signal output
rlabel metal2 s 321742 0 321798 800 6 la_data_out[83]
port 239 nsew signal output
rlabel metal2 s 325330 0 325386 800 6 la_data_out[84]
port 240 nsew signal output
rlabel metal2 s 328918 0 328974 800 6 la_data_out[85]
port 241 nsew signal output
rlabel metal2 s 332506 0 332562 800 6 la_data_out[86]
port 242 nsew signal output
rlabel metal2 s 336094 0 336150 800 6 la_data_out[87]
port 243 nsew signal output
rlabel metal2 s 339682 0 339738 800 6 la_data_out[88]
port 244 nsew signal output
rlabel metal2 s 343270 0 343326 800 6 la_data_out[89]
port 245 nsew signal output
rlabel metal2 s 52642 0 52698 800 6 la_data_out[8]
port 246 nsew signal output
rlabel metal2 s 346858 0 346914 800 6 la_data_out[90]
port 247 nsew signal output
rlabel metal2 s 350446 0 350502 800 6 la_data_out[91]
port 248 nsew signal output
rlabel metal2 s 354034 0 354090 800 6 la_data_out[92]
port 249 nsew signal output
rlabel metal2 s 357622 0 357678 800 6 la_data_out[93]
port 250 nsew signal output
rlabel metal2 s 361210 0 361266 800 6 la_data_out[94]
port 251 nsew signal output
rlabel metal2 s 364798 0 364854 800 6 la_data_out[95]
port 252 nsew signal output
rlabel metal2 s 368386 0 368442 800 6 la_data_out[96]
port 253 nsew signal output
rlabel metal2 s 371974 0 372030 800 6 la_data_out[97]
port 254 nsew signal output
rlabel metal2 s 375562 0 375618 800 6 la_data_out[98]
port 255 nsew signal output
rlabel metal2 s 379150 0 379206 800 6 la_data_out[99]
port 256 nsew signal output
rlabel metal2 s 56230 0 56286 800 6 la_data_out[9]
port 257 nsew signal output
rlabel metal2 s 25134 0 25190 800 6 la_oenb[0]
port 258 nsew signal input
rlabel metal2 s 383934 0 383990 800 6 la_oenb[100]
port 259 nsew signal input
rlabel metal2 s 387522 0 387578 800 6 la_oenb[101]
port 260 nsew signal input
rlabel metal2 s 391110 0 391166 800 6 la_oenb[102]
port 261 nsew signal input
rlabel metal2 s 394698 0 394754 800 6 la_oenb[103]
port 262 nsew signal input
rlabel metal2 s 398286 0 398342 800 6 la_oenb[104]
port 263 nsew signal input
rlabel metal2 s 401874 0 401930 800 6 la_oenb[105]
port 264 nsew signal input
rlabel metal2 s 405462 0 405518 800 6 la_oenb[106]
port 265 nsew signal input
rlabel metal2 s 409050 0 409106 800 6 la_oenb[107]
port 266 nsew signal input
rlabel metal2 s 412638 0 412694 800 6 la_oenb[108]
port 267 nsew signal input
rlabel metal2 s 416226 0 416282 800 6 la_oenb[109]
port 268 nsew signal input
rlabel metal2 s 61014 0 61070 800 6 la_oenb[10]
port 269 nsew signal input
rlabel metal2 s 419814 0 419870 800 6 la_oenb[110]
port 270 nsew signal input
rlabel metal2 s 423402 0 423458 800 6 la_oenb[111]
port 271 nsew signal input
rlabel metal2 s 426990 0 427046 800 6 la_oenb[112]
port 272 nsew signal input
rlabel metal2 s 430578 0 430634 800 6 la_oenb[113]
port 273 nsew signal input
rlabel metal2 s 434166 0 434222 800 6 la_oenb[114]
port 274 nsew signal input
rlabel metal2 s 437754 0 437810 800 6 la_oenb[115]
port 275 nsew signal input
rlabel metal2 s 441342 0 441398 800 6 la_oenb[116]
port 276 nsew signal input
rlabel metal2 s 444930 0 444986 800 6 la_oenb[117]
port 277 nsew signal input
rlabel metal2 s 448518 0 448574 800 6 la_oenb[118]
port 278 nsew signal input
rlabel metal2 s 452106 0 452162 800 6 la_oenb[119]
port 279 nsew signal input
rlabel metal2 s 64602 0 64658 800 6 la_oenb[11]
port 280 nsew signal input
rlabel metal2 s 455694 0 455750 800 6 la_oenb[120]
port 281 nsew signal input
rlabel metal2 s 459282 0 459338 800 6 la_oenb[121]
port 282 nsew signal input
rlabel metal2 s 462870 0 462926 800 6 la_oenb[122]
port 283 nsew signal input
rlabel metal2 s 466458 0 466514 800 6 la_oenb[123]
port 284 nsew signal input
rlabel metal2 s 470046 0 470102 800 6 la_oenb[124]
port 285 nsew signal input
rlabel metal2 s 473634 0 473690 800 6 la_oenb[125]
port 286 nsew signal input
rlabel metal2 s 477222 0 477278 800 6 la_oenb[126]
port 287 nsew signal input
rlabel metal2 s 480810 0 480866 800 6 la_oenb[127]
port 288 nsew signal input
rlabel metal2 s 68190 0 68246 800 6 la_oenb[12]
port 289 nsew signal input
rlabel metal2 s 71778 0 71834 800 6 la_oenb[13]
port 290 nsew signal input
rlabel metal2 s 75366 0 75422 800 6 la_oenb[14]
port 291 nsew signal input
rlabel metal2 s 78954 0 79010 800 6 la_oenb[15]
port 292 nsew signal input
rlabel metal2 s 82542 0 82598 800 6 la_oenb[16]
port 293 nsew signal input
rlabel metal2 s 86130 0 86186 800 6 la_oenb[17]
port 294 nsew signal input
rlabel metal2 s 89718 0 89774 800 6 la_oenb[18]
port 295 nsew signal input
rlabel metal2 s 93306 0 93362 800 6 la_oenb[19]
port 296 nsew signal input
rlabel metal2 s 28722 0 28778 800 6 la_oenb[1]
port 297 nsew signal input
rlabel metal2 s 96894 0 96950 800 6 la_oenb[20]
port 298 nsew signal input
rlabel metal2 s 100482 0 100538 800 6 la_oenb[21]
port 299 nsew signal input
rlabel metal2 s 104070 0 104126 800 6 la_oenb[22]
port 300 nsew signal input
rlabel metal2 s 107658 0 107714 800 6 la_oenb[23]
port 301 nsew signal input
rlabel metal2 s 111246 0 111302 800 6 la_oenb[24]
port 302 nsew signal input
rlabel metal2 s 114834 0 114890 800 6 la_oenb[25]
port 303 nsew signal input
rlabel metal2 s 118422 0 118478 800 6 la_oenb[26]
port 304 nsew signal input
rlabel metal2 s 122010 0 122066 800 6 la_oenb[27]
port 305 nsew signal input
rlabel metal2 s 125598 0 125654 800 6 la_oenb[28]
port 306 nsew signal input
rlabel metal2 s 129186 0 129242 800 6 la_oenb[29]
port 307 nsew signal input
rlabel metal2 s 32310 0 32366 800 6 la_oenb[2]
port 308 nsew signal input
rlabel metal2 s 132774 0 132830 800 6 la_oenb[30]
port 309 nsew signal input
rlabel metal2 s 136362 0 136418 800 6 la_oenb[31]
port 310 nsew signal input
rlabel metal2 s 139950 0 140006 800 6 la_oenb[32]
port 311 nsew signal input
rlabel metal2 s 143538 0 143594 800 6 la_oenb[33]
port 312 nsew signal input
rlabel metal2 s 147126 0 147182 800 6 la_oenb[34]
port 313 nsew signal input
rlabel metal2 s 150714 0 150770 800 6 la_oenb[35]
port 314 nsew signal input
rlabel metal2 s 154302 0 154358 800 6 la_oenb[36]
port 315 nsew signal input
rlabel metal2 s 157890 0 157946 800 6 la_oenb[37]
port 316 nsew signal input
rlabel metal2 s 161478 0 161534 800 6 la_oenb[38]
port 317 nsew signal input
rlabel metal2 s 165066 0 165122 800 6 la_oenb[39]
port 318 nsew signal input
rlabel metal2 s 35898 0 35954 800 6 la_oenb[3]
port 319 nsew signal input
rlabel metal2 s 168654 0 168710 800 6 la_oenb[40]
port 320 nsew signal input
rlabel metal2 s 172242 0 172298 800 6 la_oenb[41]
port 321 nsew signal input
rlabel metal2 s 175830 0 175886 800 6 la_oenb[42]
port 322 nsew signal input
rlabel metal2 s 179418 0 179474 800 6 la_oenb[43]
port 323 nsew signal input
rlabel metal2 s 183006 0 183062 800 6 la_oenb[44]
port 324 nsew signal input
rlabel metal2 s 186594 0 186650 800 6 la_oenb[45]
port 325 nsew signal input
rlabel metal2 s 190182 0 190238 800 6 la_oenb[46]
port 326 nsew signal input
rlabel metal2 s 193770 0 193826 800 6 la_oenb[47]
port 327 nsew signal input
rlabel metal2 s 197358 0 197414 800 6 la_oenb[48]
port 328 nsew signal input
rlabel metal2 s 200946 0 201002 800 6 la_oenb[49]
port 329 nsew signal input
rlabel metal2 s 39486 0 39542 800 6 la_oenb[4]
port 330 nsew signal input
rlabel metal2 s 204534 0 204590 800 6 la_oenb[50]
port 331 nsew signal input
rlabel metal2 s 208122 0 208178 800 6 la_oenb[51]
port 332 nsew signal input
rlabel metal2 s 211710 0 211766 800 6 la_oenb[52]
port 333 nsew signal input
rlabel metal2 s 215298 0 215354 800 6 la_oenb[53]
port 334 nsew signal input
rlabel metal2 s 218886 0 218942 800 6 la_oenb[54]
port 335 nsew signal input
rlabel metal2 s 222474 0 222530 800 6 la_oenb[55]
port 336 nsew signal input
rlabel metal2 s 226062 0 226118 800 6 la_oenb[56]
port 337 nsew signal input
rlabel metal2 s 229650 0 229706 800 6 la_oenb[57]
port 338 nsew signal input
rlabel metal2 s 233238 0 233294 800 6 la_oenb[58]
port 339 nsew signal input
rlabel metal2 s 236826 0 236882 800 6 la_oenb[59]
port 340 nsew signal input
rlabel metal2 s 43074 0 43130 800 6 la_oenb[5]
port 341 nsew signal input
rlabel metal2 s 240414 0 240470 800 6 la_oenb[60]
port 342 nsew signal input
rlabel metal2 s 244002 0 244058 800 6 la_oenb[61]
port 343 nsew signal input
rlabel metal2 s 247590 0 247646 800 6 la_oenb[62]
port 344 nsew signal input
rlabel metal2 s 251178 0 251234 800 6 la_oenb[63]
port 345 nsew signal input
rlabel metal2 s 254766 0 254822 800 6 la_oenb[64]
port 346 nsew signal input
rlabel metal2 s 258354 0 258410 800 6 la_oenb[65]
port 347 nsew signal input
rlabel metal2 s 261942 0 261998 800 6 la_oenb[66]
port 348 nsew signal input
rlabel metal2 s 265530 0 265586 800 6 la_oenb[67]
port 349 nsew signal input
rlabel metal2 s 269118 0 269174 800 6 la_oenb[68]
port 350 nsew signal input
rlabel metal2 s 272706 0 272762 800 6 la_oenb[69]
port 351 nsew signal input
rlabel metal2 s 46662 0 46718 800 6 la_oenb[6]
port 352 nsew signal input
rlabel metal2 s 276294 0 276350 800 6 la_oenb[70]
port 353 nsew signal input
rlabel metal2 s 279882 0 279938 800 6 la_oenb[71]
port 354 nsew signal input
rlabel metal2 s 283470 0 283526 800 6 la_oenb[72]
port 355 nsew signal input
rlabel metal2 s 287058 0 287114 800 6 la_oenb[73]
port 356 nsew signal input
rlabel metal2 s 290646 0 290702 800 6 la_oenb[74]
port 357 nsew signal input
rlabel metal2 s 294234 0 294290 800 6 la_oenb[75]
port 358 nsew signal input
rlabel metal2 s 297822 0 297878 800 6 la_oenb[76]
port 359 nsew signal input
rlabel metal2 s 301410 0 301466 800 6 la_oenb[77]
port 360 nsew signal input
rlabel metal2 s 304998 0 305054 800 6 la_oenb[78]
port 361 nsew signal input
rlabel metal2 s 308586 0 308642 800 6 la_oenb[79]
port 362 nsew signal input
rlabel metal2 s 50250 0 50306 800 6 la_oenb[7]
port 363 nsew signal input
rlabel metal2 s 312174 0 312230 800 6 la_oenb[80]
port 364 nsew signal input
rlabel metal2 s 315762 0 315818 800 6 la_oenb[81]
port 365 nsew signal input
rlabel metal2 s 319350 0 319406 800 6 la_oenb[82]
port 366 nsew signal input
rlabel metal2 s 322938 0 322994 800 6 la_oenb[83]
port 367 nsew signal input
rlabel metal2 s 326526 0 326582 800 6 la_oenb[84]
port 368 nsew signal input
rlabel metal2 s 330114 0 330170 800 6 la_oenb[85]
port 369 nsew signal input
rlabel metal2 s 333702 0 333758 800 6 la_oenb[86]
port 370 nsew signal input
rlabel metal2 s 337290 0 337346 800 6 la_oenb[87]
port 371 nsew signal input
rlabel metal2 s 340878 0 340934 800 6 la_oenb[88]
port 372 nsew signal input
rlabel metal2 s 344466 0 344522 800 6 la_oenb[89]
port 373 nsew signal input
rlabel metal2 s 53838 0 53894 800 6 la_oenb[8]
port 374 nsew signal input
rlabel metal2 s 348054 0 348110 800 6 la_oenb[90]
port 375 nsew signal input
rlabel metal2 s 351642 0 351698 800 6 la_oenb[91]
port 376 nsew signal input
rlabel metal2 s 355230 0 355286 800 6 la_oenb[92]
port 377 nsew signal input
rlabel metal2 s 358818 0 358874 800 6 la_oenb[93]
port 378 nsew signal input
rlabel metal2 s 362406 0 362462 800 6 la_oenb[94]
port 379 nsew signal input
rlabel metal2 s 365994 0 366050 800 6 la_oenb[95]
port 380 nsew signal input
rlabel metal2 s 369582 0 369638 800 6 la_oenb[96]
port 381 nsew signal input
rlabel metal2 s 373170 0 373226 800 6 la_oenb[97]
port 382 nsew signal input
rlabel metal2 s 376758 0 376814 800 6 la_oenb[98]
port 383 nsew signal input
rlabel metal2 s 380346 0 380402 800 6 la_oenb[99]
port 384 nsew signal input
rlabel metal2 s 57426 0 57482 800 6 la_oenb[9]
port 385 nsew signal input
rlabel metal4 s 4208 2128 4528 349840 6 vccd1
port 386 nsew power bidirectional
rlabel metal4 s 34928 2128 35248 349840 6 vccd1
port 386 nsew power bidirectional
rlabel metal4 s 65648 2128 65968 349840 6 vccd1
port 386 nsew power bidirectional
rlabel metal4 s 96368 2128 96688 349840 6 vccd1
port 386 nsew power bidirectional
rlabel metal4 s 127088 2128 127408 349840 6 vccd1
port 386 nsew power bidirectional
rlabel metal4 s 157808 2128 158128 349840 6 vccd1
port 386 nsew power bidirectional
rlabel metal4 s 188528 2128 188848 349840 6 vccd1
port 386 nsew power bidirectional
rlabel metal4 s 219248 2128 219568 349840 6 vccd1
port 386 nsew power bidirectional
rlabel metal4 s 249968 2128 250288 349840 6 vccd1
port 386 nsew power bidirectional
rlabel metal4 s 280688 2128 281008 349840 6 vccd1
port 386 nsew power bidirectional
rlabel metal4 s 311408 2128 311728 349840 6 vccd1
port 386 nsew power bidirectional
rlabel metal4 s 342128 2128 342448 349840 6 vccd1
port 386 nsew power bidirectional
rlabel metal4 s 372848 2128 373168 349840 6 vccd1
port 386 nsew power bidirectional
rlabel metal4 s 403568 2128 403888 349840 6 vccd1
port 386 nsew power bidirectional
rlabel metal4 s 434288 2128 434608 349840 6 vccd1
port 386 nsew power bidirectional
rlabel metal4 s 465008 2128 465328 349840 6 vccd1
port 386 nsew power bidirectional
rlabel metal4 s 495728 2128 496048 349840 6 vccd1
port 386 nsew power bidirectional
rlabel metal4 s 19568 2128 19888 349840 6 vdda1
port 387 nsew power bidirectional
rlabel metal4 s 50288 2128 50608 349840 6 vdda1
port 387 nsew power bidirectional
rlabel metal4 s 81008 2128 81328 349840 6 vdda1
port 387 nsew power bidirectional
rlabel metal4 s 111728 2128 112048 349840 6 vdda1
port 387 nsew power bidirectional
rlabel metal4 s 142448 2128 142768 349840 6 vdda1
port 387 nsew power bidirectional
rlabel metal4 s 173168 2128 173488 349840 6 vdda1
port 387 nsew power bidirectional
rlabel metal4 s 203888 2128 204208 349840 6 vdda1
port 387 nsew power bidirectional
rlabel metal4 s 234608 2128 234928 349840 6 vdda1
port 387 nsew power bidirectional
rlabel metal4 s 265328 2128 265648 349840 6 vdda1
port 387 nsew power bidirectional
rlabel metal4 s 296048 2128 296368 349840 6 vdda1
port 387 nsew power bidirectional
rlabel metal4 s 326768 2128 327088 349840 6 vdda1
port 387 nsew power bidirectional
rlabel metal4 s 357488 2128 357808 349840 6 vdda1
port 387 nsew power bidirectional
rlabel metal4 s 388208 2128 388528 349840 6 vdda1
port 387 nsew power bidirectional
rlabel metal4 s 418928 2128 419248 349840 6 vdda1
port 387 nsew power bidirectional
rlabel metal4 s 449648 2128 449968 349840 6 vdda1
port 387 nsew power bidirectional
rlabel metal4 s 480368 2128 480688 349840 6 vdda1
port 387 nsew power bidirectional
rlabel metal4 s 27248 2128 27568 349840 6 vssa1
port 388 nsew ground bidirectional
rlabel metal4 s 57968 2128 58288 349840 6 vssa1
port 388 nsew ground bidirectional
rlabel metal4 s 88688 2128 89008 349840 6 vssa1
port 388 nsew ground bidirectional
rlabel metal4 s 119408 2128 119728 349840 6 vssa1
port 388 nsew ground bidirectional
rlabel metal4 s 150128 2128 150448 349840 6 vssa1
port 388 nsew ground bidirectional
rlabel metal4 s 180848 2128 181168 349840 6 vssa1
port 388 nsew ground bidirectional
rlabel metal4 s 211568 2128 211888 349840 6 vssa1
port 388 nsew ground bidirectional
rlabel metal4 s 242288 2128 242608 349840 6 vssa1
port 388 nsew ground bidirectional
rlabel metal4 s 273008 2128 273328 349840 6 vssa1
port 388 nsew ground bidirectional
rlabel metal4 s 303728 2128 304048 349840 6 vssa1
port 388 nsew ground bidirectional
rlabel metal4 s 334448 2128 334768 349840 6 vssa1
port 388 nsew ground bidirectional
rlabel metal4 s 365168 2128 365488 349840 6 vssa1
port 388 nsew ground bidirectional
rlabel metal4 s 395888 2128 396208 349840 6 vssa1
port 388 nsew ground bidirectional
rlabel metal4 s 426608 2128 426928 349840 6 vssa1
port 388 nsew ground bidirectional
rlabel metal4 s 457328 2128 457648 349840 6 vssa1
port 388 nsew ground bidirectional
rlabel metal4 s 488048 2128 488368 349840 6 vssa1
port 388 nsew ground bidirectional
rlabel metal4 s 11888 2128 12208 349840 6 vssd1
port 389 nsew ground bidirectional
rlabel metal4 s 42608 2128 42928 349840 6 vssd1
port 389 nsew ground bidirectional
rlabel metal4 s 73328 2128 73648 349840 6 vssd1
port 389 nsew ground bidirectional
rlabel metal4 s 104048 2128 104368 349840 6 vssd1
port 389 nsew ground bidirectional
rlabel metal4 s 134768 2128 135088 349840 6 vssd1
port 389 nsew ground bidirectional
rlabel metal4 s 165488 2128 165808 349840 6 vssd1
port 389 nsew ground bidirectional
rlabel metal4 s 196208 2128 196528 349840 6 vssd1
port 389 nsew ground bidirectional
rlabel metal4 s 226928 2128 227248 349840 6 vssd1
port 389 nsew ground bidirectional
rlabel metal4 s 257648 2128 257968 349840 6 vssd1
port 389 nsew ground bidirectional
rlabel metal4 s 288368 2128 288688 349840 6 vssd1
port 389 nsew ground bidirectional
rlabel metal4 s 319088 2128 319408 349840 6 vssd1
port 389 nsew ground bidirectional
rlabel metal4 s 349808 2128 350128 349840 6 vssd1
port 389 nsew ground bidirectional
rlabel metal4 s 380528 2128 380848 349840 6 vssd1
port 389 nsew ground bidirectional
rlabel metal4 s 411248 2128 411568 349840 6 vssd1
port 389 nsew ground bidirectional
rlabel metal4 s 441968 2128 442288 349840 6 vssd1
port 389 nsew ground bidirectional
rlabel metal4 s 472688 2128 473008 349840 6 vssd1
port 389 nsew ground bidirectional
rlabel metal2 s 17958 0 18014 800 6 wb_clk_i
port 390 nsew signal input
rlabel metal2 s 19154 0 19210 800 6 wb_rst_i
port 391 nsew signal input
rlabel metal2 s 21546 0 21602 800 6 wbs_cyc_i
port 392 nsew signal input
rlabel metal2 s 20350 0 20406 800 6 wbs_stb_i
port 393 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 500000 352000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 46344762
string GDS_FILE /home/engtech/Desktop/Openlane_v2/pulse_generator_LA_v2/openlane/user_proj_example/runs/24_04_11_15_23/results/signoff/user_proj_example.magic.gds
string GDS_START 211918
<< end >>

