magic
tech sky130A
magscale 1 2
timestamp 1711496570
<< nwell >>
rect 1066 97093 98846 97414
rect 1066 96005 98846 96571
rect 1066 94917 98846 95483
rect 1066 93829 98846 94395
rect 1066 92741 98846 93307
rect 1066 91653 98846 92219
rect 1066 90565 98846 91131
rect 1066 89477 98846 90043
rect 1066 88389 98846 88955
rect 1066 87301 98846 87867
rect 1066 86213 98846 86779
rect 1066 85125 98846 85691
rect 1066 84037 98846 84603
rect 1066 82949 98846 83515
rect 1066 81861 98846 82427
rect 1066 80773 98846 81339
rect 1066 79685 98846 80251
rect 1066 78597 98846 79163
rect 1066 77509 98846 78075
rect 1066 76421 98846 76987
rect 1066 75333 98846 75899
rect 1066 74245 98846 74811
rect 1066 73157 98846 73723
rect 1066 72069 98846 72635
rect 1066 70981 98846 71547
rect 1066 69893 98846 70459
rect 1066 68805 98846 69371
rect 1066 67717 98846 68283
rect 1066 66629 98846 67195
rect 1066 65541 98846 66107
rect 1066 64453 98846 65019
rect 1066 63365 98846 63931
rect 1066 62277 98846 62843
rect 1066 61189 98846 61755
rect 1066 60101 98846 60667
rect 1066 59013 98846 59579
rect 1066 57925 98846 58491
rect 1066 56837 98846 57403
rect 1066 55749 98846 56315
rect 1066 54661 98846 55227
rect 1066 53573 98846 54139
rect 1066 52485 98846 53051
rect 1066 51397 98846 51963
rect 1066 50309 98846 50875
rect 1066 49221 98846 49787
rect 1066 48133 98846 48699
rect 1066 47045 98846 47611
rect 1066 45957 98846 46523
rect 1066 44869 98846 45435
rect 1066 43781 98846 44347
rect 1066 42693 98846 43259
rect 1066 41605 98846 42171
rect 1066 40517 98846 41083
rect 1066 39429 98846 39995
rect 1066 38341 98846 38907
rect 1066 37253 98846 37819
rect 1066 36165 98846 36731
rect 1066 35077 98846 35643
rect 1066 33989 98846 34555
rect 1066 32901 98846 33467
rect 1066 31813 98846 32379
rect 1066 30725 98846 31291
rect 1066 29637 98846 30203
rect 1066 28549 98846 29115
rect 1066 27461 98846 28027
rect 1066 26373 98846 26939
rect 1066 25285 98846 25851
rect 1066 24197 98846 24763
rect 1066 23109 98846 23675
rect 1066 22021 98846 22587
rect 1066 20933 98846 21499
rect 1066 19845 98846 20411
rect 1066 18757 98846 19323
rect 1066 17669 98846 18235
rect 1066 16581 98846 17147
rect 1066 15493 98846 16059
rect 1066 14405 98846 14971
rect 1066 13317 98846 13883
rect 1066 12229 98846 12795
rect 1066 11141 98846 11707
rect 1066 10053 98846 10619
rect 1066 8965 98846 9531
rect 1066 7877 98846 8443
rect 1066 6789 98846 7355
rect 1066 5701 98846 6267
rect 1066 4613 98846 5179
rect 1066 3525 98846 4091
rect 1066 2437 98846 3003
<< obsli1 >>
rect 1104 2159 98808 97393
<< obsm1 >>
rect 1104 1640 98808 97424
<< metal2 >>
rect 3698 0 3754 800
rect 9862 0 9918 800
rect 16026 0 16082 800
rect 22190 0 22246 800
rect 28354 0 28410 800
rect 34518 0 34574 800
rect 40682 0 40738 800
rect 46846 0 46902 800
rect 53010 0 53066 800
rect 59174 0 59230 800
rect 65338 0 65394 800
rect 71502 0 71558 800
rect 77666 0 77722 800
rect 83830 0 83886 800
rect 89994 0 90050 800
rect 96158 0 96214 800
<< obsm2 >>
rect 3698 856 96682 97413
rect 3810 800 9806 856
rect 9974 800 15970 856
rect 16138 800 22134 856
rect 22302 800 28298 856
rect 28466 800 34462 856
rect 34630 800 40626 856
rect 40794 800 46790 856
rect 46958 800 52954 856
rect 53122 800 59118 856
rect 59286 800 65282 856
rect 65450 800 71446 856
rect 71614 800 77610 856
rect 77778 800 83774 856
rect 83942 800 89938 856
rect 90106 800 96102 856
rect 96270 800 96682 856
<< obsm3 >>
rect 3693 2143 96686 97409
<< metal4 >>
rect 4208 2128 4528 97424
rect 19568 2128 19888 97424
rect 34928 2128 35248 97424
rect 50288 2128 50608 97424
rect 65648 2128 65968 97424
rect 81008 2128 81328 97424
rect 96368 2128 96688 97424
<< labels >>
rlabel metal2 s 34518 0 34574 800 6 la_data_in[0]
port 1 nsew signal input
rlabel metal2 s 46846 0 46902 800 6 la_data_in[1]
port 2 nsew signal input
rlabel metal2 s 59174 0 59230 800 6 la_data_in[2]
port 3 nsew signal input
rlabel metal2 s 71502 0 71558 800 6 la_data_in[3]
port 4 nsew signal input
rlabel metal2 s 83830 0 83886 800 6 la_data_in[4]
port 5 nsew signal input
rlabel metal2 s 28354 0 28410 800 6 la_data_out
port 6 nsew signal output
rlabel metal2 s 40682 0 40738 800 6 la_oenb[0]
port 7 nsew signal input
rlabel metal2 s 53010 0 53066 800 6 la_oenb[1]
port 8 nsew signal input
rlabel metal2 s 65338 0 65394 800 6 la_oenb[2]
port 9 nsew signal input
rlabel metal2 s 77666 0 77722 800 6 la_oenb[3]
port 10 nsew signal input
rlabel metal2 s 89994 0 90050 800 6 la_oenb[4]
port 11 nsew signal input
rlabel metal2 s 96158 0 96214 800 6 la_oenb[5]
port 12 nsew signal input
rlabel metal4 s 4208 2128 4528 97424 6 vccd1
port 13 nsew power bidirectional
rlabel metal4 s 34928 2128 35248 97424 6 vccd1
port 13 nsew power bidirectional
rlabel metal4 s 65648 2128 65968 97424 6 vccd1
port 13 nsew power bidirectional
rlabel metal4 s 96368 2128 96688 97424 6 vccd1
port 13 nsew power bidirectional
rlabel metal4 s 19568 2128 19888 97424 6 vssd1
port 14 nsew ground bidirectional
rlabel metal4 s 50288 2128 50608 97424 6 vssd1
port 14 nsew ground bidirectional
rlabel metal4 s 81008 2128 81328 97424 6 vssd1
port 14 nsew ground bidirectional
rlabel metal2 s 3698 0 3754 800 6 wb_clk_i
port 15 nsew signal input
rlabel metal2 s 9862 0 9918 800 6 wb_rst_i
port 16 nsew signal input
rlabel metal2 s 16026 0 16082 800 6 wbs_cyc_i
port 17 nsew signal input
rlabel metal2 s 22190 0 22246 800 6 wbs_stb_i
port 18 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 100000 100000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 2871316
string GDS_FILE /home/engtech/Desktop/Openlane_v2/pulse_generator_LA/openlane/user_proj_example/runs/24_03_26_18_41/results/signoff/user_proj_example.magic.gds
string GDS_START 201568
<< end >>

