VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO user_proj_example
  CLASS BLOCK ;
  FOREIGN user_proj_example ;
  ORIGIN 0.000 0.000 ;
  SIZE 500.000 BY 500.000 ;
  PIN la_data_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 172.590 0.000 172.870 4.000 ;
    END
  END la_data_in[0]
  PIN la_data_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 234.230 0.000 234.510 4.000 ;
    END
  END la_data_in[1]
  PIN la_data_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 295.870 0.000 296.150 4.000 ;
    END
  END la_data_in[2]
  PIN la_data_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 357.510 0.000 357.790 4.000 ;
    END
  END la_data_in[3]
  PIN la_data_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 419.150 0.000 419.430 4.000 ;
    END
  END la_data_in[4]
  PIN la_data_out
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 141.770 0.000 142.050 4.000 ;
    END
  END la_data_out
  PIN la_oenb[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 203.410 0.000 203.690 4.000 ;
    END
  END la_oenb[0]
  PIN la_oenb[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 265.050 0.000 265.330 4.000 ;
    END
  END la_oenb[1]
  PIN la_oenb[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 326.690 0.000 326.970 4.000 ;
    END
  END la_oenb[2]
  PIN la_oenb[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 388.330 0.000 388.610 4.000 ;
    END
  END la_oenb[3]
  PIN la_oenb[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 449.970 0.000 450.250 4.000 ;
    END
  END la_oenb[4]
  PIN la_oenb[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 480.790 0.000 481.070 4.000 ;
    END
  END la_oenb[5]
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 487.120 ;
    END
    PORT
      LAYER met4 ;
        RECT 174.640 10.640 176.240 487.120 ;
    END
    PORT
      LAYER met4 ;
        RECT 328.240 10.640 329.840 487.120 ;
    END
    PORT
      LAYER met4 ;
        RECT 481.840 10.640 483.440 487.120 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 97.840 10.640 99.440 487.120 ;
    END
    PORT
      LAYER met4 ;
        RECT 251.440 10.640 253.040 487.120 ;
    END
    PORT
      LAYER met4 ;
        RECT 405.040 10.640 406.640 487.120 ;
    END
  END vssd1
  PIN wb_clk_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 2.173500 ;
    PORT
      LAYER met2 ;
        RECT 18.490 0.000 18.770 4.000 ;
    END
  END wb_clk_i
  PIN wb_rst_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 49.310 0.000 49.590 4.000 ;
    END
  END wb_rst_i
  PIN wbs_cyc_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 80.130 0.000 80.410 4.000 ;
    END
  END wbs_cyc_i
  PIN wbs_stb_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 110.950 0.000 111.230 4.000 ;
    END
  END wbs_stb_i
  OBS
      LAYER nwell ;
        RECT 5.330 485.465 494.230 487.070 ;
        RECT 5.330 480.025 494.230 482.855 ;
        RECT 5.330 474.585 494.230 477.415 ;
        RECT 5.330 469.145 494.230 471.975 ;
        RECT 5.330 463.705 494.230 466.535 ;
        RECT 5.330 458.265 494.230 461.095 ;
        RECT 5.330 452.825 494.230 455.655 ;
        RECT 5.330 447.385 494.230 450.215 ;
        RECT 5.330 441.945 494.230 444.775 ;
        RECT 5.330 436.505 494.230 439.335 ;
        RECT 5.330 431.065 494.230 433.895 ;
        RECT 5.330 425.625 494.230 428.455 ;
        RECT 5.330 420.185 494.230 423.015 ;
        RECT 5.330 414.745 494.230 417.575 ;
        RECT 5.330 409.305 494.230 412.135 ;
        RECT 5.330 403.865 494.230 406.695 ;
        RECT 5.330 398.425 494.230 401.255 ;
        RECT 5.330 392.985 494.230 395.815 ;
        RECT 5.330 387.545 494.230 390.375 ;
        RECT 5.330 382.105 494.230 384.935 ;
        RECT 5.330 376.665 494.230 379.495 ;
        RECT 5.330 371.225 494.230 374.055 ;
        RECT 5.330 365.785 494.230 368.615 ;
        RECT 5.330 360.345 494.230 363.175 ;
        RECT 5.330 354.905 494.230 357.735 ;
        RECT 5.330 349.465 494.230 352.295 ;
        RECT 5.330 344.025 494.230 346.855 ;
        RECT 5.330 338.585 494.230 341.415 ;
        RECT 5.330 333.145 494.230 335.975 ;
        RECT 5.330 327.705 494.230 330.535 ;
        RECT 5.330 322.265 494.230 325.095 ;
        RECT 5.330 316.825 494.230 319.655 ;
        RECT 5.330 311.385 494.230 314.215 ;
        RECT 5.330 305.945 494.230 308.775 ;
        RECT 5.330 300.505 494.230 303.335 ;
        RECT 5.330 295.065 494.230 297.895 ;
        RECT 5.330 289.625 494.230 292.455 ;
        RECT 5.330 284.185 494.230 287.015 ;
        RECT 5.330 278.745 494.230 281.575 ;
        RECT 5.330 273.305 494.230 276.135 ;
        RECT 5.330 267.865 494.230 270.695 ;
        RECT 5.330 262.425 494.230 265.255 ;
        RECT 5.330 256.985 494.230 259.815 ;
        RECT 5.330 251.545 494.230 254.375 ;
        RECT 5.330 246.105 494.230 248.935 ;
        RECT 5.330 240.665 494.230 243.495 ;
        RECT 5.330 235.225 494.230 238.055 ;
        RECT 5.330 229.785 494.230 232.615 ;
        RECT 5.330 224.345 494.230 227.175 ;
        RECT 5.330 218.905 494.230 221.735 ;
        RECT 5.330 213.465 494.230 216.295 ;
        RECT 5.330 208.025 494.230 210.855 ;
        RECT 5.330 202.585 494.230 205.415 ;
        RECT 5.330 197.145 494.230 199.975 ;
        RECT 5.330 191.705 494.230 194.535 ;
        RECT 5.330 186.265 494.230 189.095 ;
        RECT 5.330 180.825 494.230 183.655 ;
        RECT 5.330 175.385 494.230 178.215 ;
        RECT 5.330 169.945 494.230 172.775 ;
        RECT 5.330 164.505 494.230 167.335 ;
        RECT 5.330 159.065 494.230 161.895 ;
        RECT 5.330 153.625 494.230 156.455 ;
        RECT 5.330 148.185 494.230 151.015 ;
        RECT 5.330 142.745 494.230 145.575 ;
        RECT 5.330 137.305 494.230 140.135 ;
        RECT 5.330 131.865 494.230 134.695 ;
        RECT 5.330 126.425 494.230 129.255 ;
        RECT 5.330 120.985 494.230 123.815 ;
        RECT 5.330 115.545 494.230 118.375 ;
        RECT 5.330 110.105 494.230 112.935 ;
        RECT 5.330 104.665 494.230 107.495 ;
        RECT 5.330 99.225 494.230 102.055 ;
        RECT 5.330 93.785 494.230 96.615 ;
        RECT 5.330 88.345 494.230 91.175 ;
        RECT 5.330 82.905 494.230 85.735 ;
        RECT 5.330 77.465 494.230 80.295 ;
        RECT 5.330 72.025 494.230 74.855 ;
        RECT 5.330 66.585 494.230 69.415 ;
        RECT 5.330 61.145 494.230 63.975 ;
        RECT 5.330 55.705 494.230 58.535 ;
        RECT 5.330 50.265 494.230 53.095 ;
        RECT 5.330 44.825 494.230 47.655 ;
        RECT 5.330 39.385 494.230 42.215 ;
        RECT 5.330 33.945 494.230 36.775 ;
        RECT 5.330 28.505 494.230 31.335 ;
        RECT 5.330 23.065 494.230 25.895 ;
        RECT 5.330 17.625 494.230 20.455 ;
        RECT 5.330 12.185 494.230 15.015 ;
      LAYER li1 ;
        RECT 5.520 10.795 494.040 486.965 ;
      LAYER met1 ;
        RECT 5.520 8.200 494.040 487.120 ;
      LAYER met2 ;
        RECT 18.490 4.280 483.410 487.065 ;
        RECT 19.050 4.000 49.030 4.280 ;
        RECT 49.870 4.000 79.850 4.280 ;
        RECT 80.690 4.000 110.670 4.280 ;
        RECT 111.510 4.000 141.490 4.280 ;
        RECT 142.330 4.000 172.310 4.280 ;
        RECT 173.150 4.000 203.130 4.280 ;
        RECT 203.970 4.000 233.950 4.280 ;
        RECT 234.790 4.000 264.770 4.280 ;
        RECT 265.610 4.000 295.590 4.280 ;
        RECT 296.430 4.000 326.410 4.280 ;
        RECT 327.250 4.000 357.230 4.280 ;
        RECT 358.070 4.000 388.050 4.280 ;
        RECT 388.890 4.000 418.870 4.280 ;
        RECT 419.710 4.000 449.690 4.280 ;
        RECT 450.530 4.000 480.510 4.280 ;
        RECT 481.350 4.000 483.410 4.280 ;
      LAYER met3 ;
        RECT 18.465 10.715 483.430 487.045 ;
  END
END user_proj_example
END LIBRARY

